// This  Verilog HDL  source  file was  automatically generated
// by C++ model based on VPP library. Modification of this file
// is possible, but if you want to keep it in sync with the C++
// model,  please  modify  the model and re-generate this file.
// VPP library web-page: http://www.phys.ufl.edu/~madorsky/vpp/

// Author    : ise
// File name : collider.v
// Timestamp : Fri Sep 10 20:09:53 2021

module collider
(
    qp0,
    qp1,
    qp2,
    qp3,
    w1,
    w2,
    q1,
    q2,
    v1,
    v2,
    clk
);

    input [111:0] qp0;
    input [111:0] qp1;
    input [111:0] qp2;
    input [111:0] qp3;
    output [6:0] w1;
    reg    [6:0] w1;
    output [6:0] w2;
    reg    [6:0] w2;
    output [1:0] q1;
    reg    [1:0] q1;
    output [1:0] q2;
    reg    [1:0] q2;
    output v1;
    reg    v1;
    output v2;
    reg    v2;
    input clk;

    reg [6:0] n3_1;
    reg [6:0] n3_2;
    reg [6:0] n2_1;
    reg [6:0] n2_2;
    reg [6:0] n1_1;
    reg [6:0] n1_2;
    reg [6:0] n0_1;
    reg [6:0] n0_2;
    always @(qp0 or qp1 or qp2 or qp3) 
    begin
        n3_1 = 7'h7f;
        n2_1 = 7'h7f;
        n1_1 = 7'h7f;
        n0_1 = 7'h7f;
        if (qp3[0]) n3_1 = 0;
        if (qp2[0]) n2_1 = 0;
        if (qp1[0]) n1_1 = 0;
        if (qp0[0]) n0_1 = 0;
        if (qp3[1]) n3_1 = 1;
        if (qp2[1]) n2_1 = 1;
        if (qp1[1]) n1_1 = 1;
        if (qp0[1]) n0_1 = 1;
        if (qp3[2]) n3_1 = 2;
        if (qp2[2]) n2_1 = 2;
        if (qp1[2]) n1_1 = 2;
        if (qp0[2]) n0_1 = 2;
        if (qp3[3]) n3_1 = 3;
        if (qp2[3]) n2_1 = 3;
        if (qp1[3]) n1_1 = 3;
        if (qp0[3]) n0_1 = 3;
        if (qp3[4]) n3_1 = 4;
        if (qp2[4]) n2_1 = 4;
        if (qp1[4]) n1_1 = 4;
        if (qp0[4]) n0_1 = 4;
        if (qp3[5]) n3_1 = 5;
        if (qp2[5]) n2_1 = 5;
        if (qp1[5]) n1_1 = 5;
        if (qp0[5]) n0_1 = 5;
        if (qp3[6]) n3_1 = 6;
        if (qp2[6]) n2_1 = 6;
        if (qp1[6]) n1_1 = 6;
        if (qp0[6]) n0_1 = 6;
        if (qp3[7]) n3_1 = 7;
        if (qp2[7]) n2_1 = 7;
        if (qp1[7]) n1_1 = 7;
        if (qp0[7]) n0_1 = 7;
        if (qp3[8]) n3_1 = 8;
        if (qp2[8]) n2_1 = 8;
        if (qp1[8]) n1_1 = 8;
        if (qp0[8]) n0_1 = 8;
        if (qp3[9]) n3_1 = 9;
        if (qp2[9]) n2_1 = 9;
        if (qp1[9]) n1_1 = 9;
        if (qp0[9]) n0_1 = 9;
        if (qp3[10]) n3_1 = 10;
        if (qp2[10]) n2_1 = 10;
        if (qp1[10]) n1_1 = 10;
        if (qp0[10]) n0_1 = 10;
        if (qp3[11]) n3_1 = 11;
        if (qp2[11]) n2_1 = 11;
        if (qp1[11]) n1_1 = 11;
        if (qp0[11]) n0_1 = 11;
        if (qp3[12]) n3_1 = 12;
        if (qp2[12]) n2_1 = 12;
        if (qp1[12]) n1_1 = 12;
        if (qp0[12]) n0_1 = 12;
        if (qp3[13]) n3_1 = 13;
        if (qp2[13]) n2_1 = 13;
        if (qp1[13]) n1_1 = 13;
        if (qp0[13]) n0_1 = 13;
        if (qp3[14]) n3_1 = 14;
        if (qp2[14]) n2_1 = 14;
        if (qp1[14]) n1_1 = 14;
        if (qp0[14]) n0_1 = 14;
        if (qp3[15]) n3_1 = 15;
        if (qp2[15]) n2_1 = 15;
        if (qp1[15]) n1_1 = 15;
        if (qp0[15]) n0_1 = 15;
        if (qp3[16]) n3_1 = 16;
        if (qp2[16]) n2_1 = 16;
        if (qp1[16]) n1_1 = 16;
        if (qp0[16]) n0_1 = 16;
        if (qp3[17]) n3_1 = 17;
        if (qp2[17]) n2_1 = 17;
        if (qp1[17]) n1_1 = 17;
        if (qp0[17]) n0_1 = 17;
        if (qp3[18]) n3_1 = 18;
        if (qp2[18]) n2_1 = 18;
        if (qp1[18]) n1_1 = 18;
        if (qp0[18]) n0_1 = 18;
        if (qp3[19]) n3_1 = 19;
        if (qp2[19]) n2_1 = 19;
        if (qp1[19]) n1_1 = 19;
        if (qp0[19]) n0_1 = 19;
        if (qp3[20]) n3_1 = 20;
        if (qp2[20]) n2_1 = 20;
        if (qp1[20]) n1_1 = 20;
        if (qp0[20]) n0_1 = 20;
        if (qp3[21]) n3_1 = 21;
        if (qp2[21]) n2_1 = 21;
        if (qp1[21]) n1_1 = 21;
        if (qp0[21]) n0_1 = 21;
        if (qp3[22]) n3_1 = 22;
        if (qp2[22]) n2_1 = 22;
        if (qp1[22]) n1_1 = 22;
        if (qp0[22]) n0_1 = 22;
        if (qp3[23]) n3_1 = 23;
        if (qp2[23]) n2_1 = 23;
        if (qp1[23]) n1_1 = 23;
        if (qp0[23]) n0_1 = 23;
        if (qp3[24]) n3_1 = 24;
        if (qp2[24]) n2_1 = 24;
        if (qp1[24]) n1_1 = 24;
        if (qp0[24]) n0_1 = 24;
        if (qp3[25]) n3_1 = 25;
        if (qp2[25]) n2_1 = 25;
        if (qp1[25]) n1_1 = 25;
        if (qp0[25]) n0_1 = 25;
        if (qp3[26]) n3_1 = 26;
        if (qp2[26]) n2_1 = 26;
        if (qp1[26]) n1_1 = 26;
        if (qp0[26]) n0_1 = 26;
        if (qp3[27]) n3_1 = 27;
        if (qp2[27]) n2_1 = 27;
        if (qp1[27]) n1_1 = 27;
        if (qp0[27]) n0_1 = 27;
        if (qp3[28]) n3_1 = 28;
        if (qp2[28]) n2_1 = 28;
        if (qp1[28]) n1_1 = 28;
        if (qp0[28]) n0_1 = 28;
        if (qp3[29]) n3_1 = 29;
        if (qp2[29]) n2_1 = 29;
        if (qp1[29]) n1_1 = 29;
        if (qp0[29]) n0_1 = 29;
        if (qp3[30]) n3_1 = 30;
        if (qp2[30]) n2_1 = 30;
        if (qp1[30]) n1_1 = 30;
        if (qp0[30]) n0_1 = 30;
        if (qp3[31]) n3_1 = 31;
        if (qp2[31]) n2_1 = 31;
        if (qp1[31]) n1_1 = 31;
        if (qp0[31]) n0_1 = 31;
        if (qp3[32]) n3_1 = 32;
        if (qp2[32]) n2_1 = 32;
        if (qp1[32]) n1_1 = 32;
        if (qp0[32]) n0_1 = 32;
        if (qp3[33]) n3_1 = 33;
        if (qp2[33]) n2_1 = 33;
        if (qp1[33]) n1_1 = 33;
        if (qp0[33]) n0_1 = 33;
        if (qp3[34]) n3_1 = 34;
        if (qp2[34]) n2_1 = 34;
        if (qp1[34]) n1_1 = 34;
        if (qp0[34]) n0_1 = 34;
        if (qp3[35]) n3_1 = 35;
        if (qp2[35]) n2_1 = 35;
        if (qp1[35]) n1_1 = 35;
        if (qp0[35]) n0_1 = 35;
        if (qp3[36]) n3_1 = 36;
        if (qp2[36]) n2_1 = 36;
        if (qp1[36]) n1_1 = 36;
        if (qp0[36]) n0_1 = 36;
        if (qp3[37]) n3_1 = 37;
        if (qp2[37]) n2_1 = 37;
        if (qp1[37]) n1_1 = 37;
        if (qp0[37]) n0_1 = 37;
        if (qp3[38]) n3_1 = 38;
        if (qp2[38]) n2_1 = 38;
        if (qp1[38]) n1_1 = 38;
        if (qp0[38]) n0_1 = 38;
        if (qp3[39]) n3_1 = 39;
        if (qp2[39]) n2_1 = 39;
        if (qp1[39]) n1_1 = 39;
        if (qp0[39]) n0_1 = 39;
        if (qp3[40]) n3_1 = 40;
        if (qp2[40]) n2_1 = 40;
        if (qp1[40]) n1_1 = 40;
        if (qp0[40]) n0_1 = 40;
        if (qp3[41]) n3_1 = 41;
        if (qp2[41]) n2_1 = 41;
        if (qp1[41]) n1_1 = 41;
        if (qp0[41]) n0_1 = 41;
        if (qp3[42]) n3_1 = 42;
        if (qp2[42]) n2_1 = 42;
        if (qp1[42]) n1_1 = 42;
        if (qp0[42]) n0_1 = 42;
        if (qp3[43]) n3_1 = 43;
        if (qp2[43]) n2_1 = 43;
        if (qp1[43]) n1_1 = 43;
        if (qp0[43]) n0_1 = 43;
        if (qp3[44]) n3_1 = 44;
        if (qp2[44]) n2_1 = 44;
        if (qp1[44]) n1_1 = 44;
        if (qp0[44]) n0_1 = 44;
        if (qp3[45]) n3_1 = 45;
        if (qp2[45]) n2_1 = 45;
        if (qp1[45]) n1_1 = 45;
        if (qp0[45]) n0_1 = 45;
        if (qp3[46]) n3_1 = 46;
        if (qp2[46]) n2_1 = 46;
        if (qp1[46]) n1_1 = 46;
        if (qp0[46]) n0_1 = 46;
        if (qp3[47]) n3_1 = 47;
        if (qp2[47]) n2_1 = 47;
        if (qp1[47]) n1_1 = 47;
        if (qp0[47]) n0_1 = 47;
        if (qp3[48]) n3_1 = 48;
        if (qp2[48]) n2_1 = 48;
        if (qp1[48]) n1_1 = 48;
        if (qp0[48]) n0_1 = 48;
        if (qp3[49]) n3_1 = 49;
        if (qp2[49]) n2_1 = 49;
        if (qp1[49]) n1_1 = 49;
        if (qp0[49]) n0_1 = 49;
        if (qp3[50]) n3_1 = 50;
        if (qp2[50]) n2_1 = 50;
        if (qp1[50]) n1_1 = 50;
        if (qp0[50]) n0_1 = 50;
        if (qp3[51]) n3_1 = 51;
        if (qp2[51]) n2_1 = 51;
        if (qp1[51]) n1_1 = 51;
        if (qp0[51]) n0_1 = 51;
        if (qp3[52]) n3_1 = 52;
        if (qp2[52]) n2_1 = 52;
        if (qp1[52]) n1_1 = 52;
        if (qp0[52]) n0_1 = 52;
        if (qp3[53]) n3_1 = 53;
        if (qp2[53]) n2_1 = 53;
        if (qp1[53]) n1_1 = 53;
        if (qp0[53]) n0_1 = 53;
        if (qp3[54]) n3_1 = 54;
        if (qp2[54]) n2_1 = 54;
        if (qp1[54]) n1_1 = 54;
        if (qp0[54]) n0_1 = 54;
        if (qp3[55]) n3_1 = 55;
        if (qp2[55]) n2_1 = 55;
        if (qp1[55]) n1_1 = 55;
        if (qp0[55]) n0_1 = 55;
        if (qp3[56]) n3_1 = 56;
        if (qp2[56]) n2_1 = 56;
        if (qp1[56]) n1_1 = 56;
        if (qp0[56]) n0_1 = 56;
        if (qp3[57]) n3_1 = 57;
        if (qp2[57]) n2_1 = 57;
        if (qp1[57]) n1_1 = 57;
        if (qp0[57]) n0_1 = 57;
        if (qp3[58]) n3_1 = 58;
        if (qp2[58]) n2_1 = 58;
        if (qp1[58]) n1_1 = 58;
        if (qp0[58]) n0_1 = 58;
        if (qp3[59]) n3_1 = 59;
        if (qp2[59]) n2_1 = 59;
        if (qp1[59]) n1_1 = 59;
        if (qp0[59]) n0_1 = 59;
        if (qp3[60]) n3_1 = 60;
        if (qp2[60]) n2_1 = 60;
        if (qp1[60]) n1_1 = 60;
        if (qp0[60]) n0_1 = 60;
        if (qp3[61]) n3_1 = 61;
        if (qp2[61]) n2_1 = 61;
        if (qp1[61]) n1_1 = 61;
        if (qp0[61]) n0_1 = 61;
        if (qp3[62]) n3_1 = 62;
        if (qp2[62]) n2_1 = 62;
        if (qp1[62]) n1_1 = 62;
        if (qp0[62]) n0_1 = 62;
        if (qp3[63]) n3_1 = 63;
        if (qp2[63]) n2_1 = 63;
        if (qp1[63]) n1_1 = 63;
        if (qp0[63]) n0_1 = 63;
        if (qp3[64]) n3_1 = 64;
        if (qp2[64]) n2_1 = 64;
        if (qp1[64]) n1_1 = 64;
        if (qp0[64]) n0_1 = 64;
        if (qp3[65]) n3_1 = 65;
        if (qp2[65]) n2_1 = 65;
        if (qp1[65]) n1_1 = 65;
        if (qp0[65]) n0_1 = 65;
        if (qp3[66]) n3_1 = 66;
        if (qp2[66]) n2_1 = 66;
        if (qp1[66]) n1_1 = 66;
        if (qp0[66]) n0_1 = 66;
        if (qp3[67]) n3_1 = 67;
        if (qp2[67]) n2_1 = 67;
        if (qp1[67]) n1_1 = 67;
        if (qp0[67]) n0_1 = 67;
        if (qp3[68]) n3_1 = 68;
        if (qp2[68]) n2_1 = 68;
        if (qp1[68]) n1_1 = 68;
        if (qp0[68]) n0_1 = 68;
        if (qp3[69]) n3_1 = 69;
        if (qp2[69]) n2_1 = 69;
        if (qp1[69]) n1_1 = 69;
        if (qp0[69]) n0_1 = 69;
        if (qp3[70]) n3_1 = 70;
        if (qp2[70]) n2_1 = 70;
        if (qp1[70]) n1_1 = 70;
        if (qp0[70]) n0_1 = 70;
        if (qp3[71]) n3_1 = 71;
        if (qp2[71]) n2_1 = 71;
        if (qp1[71]) n1_1 = 71;
        if (qp0[71]) n0_1 = 71;
        if (qp3[72]) n3_1 = 72;
        if (qp2[72]) n2_1 = 72;
        if (qp1[72]) n1_1 = 72;
        if (qp0[72]) n0_1 = 72;
        if (qp3[73]) n3_1 = 73;
        if (qp2[73]) n2_1 = 73;
        if (qp1[73]) n1_1 = 73;
        if (qp0[73]) n0_1 = 73;
        if (qp3[74]) n3_1 = 74;
        if (qp2[74]) n2_1 = 74;
        if (qp1[74]) n1_1 = 74;
        if (qp0[74]) n0_1 = 74;
        if (qp3[75]) n3_1 = 75;
        if (qp2[75]) n2_1 = 75;
        if (qp1[75]) n1_1 = 75;
        if (qp0[75]) n0_1 = 75;
        if (qp3[76]) n3_1 = 76;
        if (qp2[76]) n2_1 = 76;
        if (qp1[76]) n1_1 = 76;
        if (qp0[76]) n0_1 = 76;
        if (qp3[77]) n3_1 = 77;
        if (qp2[77]) n2_1 = 77;
        if (qp1[77]) n1_1 = 77;
        if (qp0[77]) n0_1 = 77;
        if (qp3[78]) n3_1 = 78;
        if (qp2[78]) n2_1 = 78;
        if (qp1[78]) n1_1 = 78;
        if (qp0[78]) n0_1 = 78;
        if (qp3[79]) n3_1 = 79;
        if (qp2[79]) n2_1 = 79;
        if (qp1[79]) n1_1 = 79;
        if (qp0[79]) n0_1 = 79;
        if (qp3[80]) n3_1 = 80;
        if (qp2[80]) n2_1 = 80;
        if (qp1[80]) n1_1 = 80;
        if (qp0[80]) n0_1 = 80;
        if (qp3[81]) n3_1 = 81;
        if (qp2[81]) n2_1 = 81;
        if (qp1[81]) n1_1 = 81;
        if (qp0[81]) n0_1 = 81;
        if (qp3[82]) n3_1 = 82;
        if (qp2[82]) n2_1 = 82;
        if (qp1[82]) n1_1 = 82;
        if (qp0[82]) n0_1 = 82;
        if (qp3[83]) n3_1 = 83;
        if (qp2[83]) n2_1 = 83;
        if (qp1[83]) n1_1 = 83;
        if (qp0[83]) n0_1 = 83;
        if (qp3[84]) n3_1 = 84;
        if (qp2[84]) n2_1 = 84;
        if (qp1[84]) n1_1 = 84;
        if (qp0[84]) n0_1 = 84;
        if (qp3[85]) n3_1 = 85;
        if (qp2[85]) n2_1 = 85;
        if (qp1[85]) n1_1 = 85;
        if (qp0[85]) n0_1 = 85;
        if (qp3[86]) n3_1 = 86;
        if (qp2[86]) n2_1 = 86;
        if (qp1[86]) n1_1 = 86;
        if (qp0[86]) n0_1 = 86;
        if (qp3[87]) n3_1 = 87;
        if (qp2[87]) n2_1 = 87;
        if (qp1[87]) n1_1 = 87;
        if (qp0[87]) n0_1 = 87;
        if (qp3[88]) n3_1 = 88;
        if (qp2[88]) n2_1 = 88;
        if (qp1[88]) n1_1 = 88;
        if (qp0[88]) n0_1 = 88;
        if (qp3[89]) n3_1 = 89;
        if (qp2[89]) n2_1 = 89;
        if (qp1[89]) n1_1 = 89;
        if (qp0[89]) n0_1 = 89;
        if (qp3[90]) n3_1 = 90;
        if (qp2[90]) n2_1 = 90;
        if (qp1[90]) n1_1 = 90;
        if (qp0[90]) n0_1 = 90;
        if (qp3[91]) n3_1 = 91;
        if (qp2[91]) n2_1 = 91;
        if (qp1[91]) n1_1 = 91;
        if (qp0[91]) n0_1 = 91;
        if (qp3[92]) n3_1 = 92;
        if (qp2[92]) n2_1 = 92;
        if (qp1[92]) n1_1 = 92;
        if (qp0[92]) n0_1 = 92;
        if (qp3[93]) n3_1 = 93;
        if (qp2[93]) n2_1 = 93;
        if (qp1[93]) n1_1 = 93;
        if (qp0[93]) n0_1 = 93;
        if (qp3[94]) n3_1 = 94;
        if (qp2[94]) n2_1 = 94;
        if (qp1[94]) n1_1 = 94;
        if (qp0[94]) n0_1 = 94;
        if (qp3[95]) n3_1 = 95;
        if (qp2[95]) n2_1 = 95;
        if (qp1[95]) n1_1 = 95;
        if (qp0[95]) n0_1 = 95;
        if (qp3[96]) n3_1 = 96;
        if (qp2[96]) n2_1 = 96;
        if (qp1[96]) n1_1 = 96;
        if (qp0[96]) n0_1 = 96;
        if (qp3[97]) n3_1 = 97;
        if (qp2[97]) n2_1 = 97;
        if (qp1[97]) n1_1 = 97;
        if (qp0[97]) n0_1 = 97;
        if (qp3[98]) n3_1 = 98;
        if (qp2[98]) n2_1 = 98;
        if (qp1[98]) n1_1 = 98;
        if (qp0[98]) n0_1 = 98;
        if (qp3[99]) n3_1 = 99;
        if (qp2[99]) n2_1 = 99;
        if (qp1[99]) n1_1 = 99;
        if (qp0[99]) n0_1 = 99;
        if (qp3[100]) n3_1 = 100;
        if (qp2[100]) n2_1 = 100;
        if (qp1[100]) n1_1 = 100;
        if (qp0[100]) n0_1 = 100;
        if (qp3[101]) n3_1 = 101;
        if (qp2[101]) n2_1 = 101;
        if (qp1[101]) n1_1 = 101;
        if (qp0[101]) n0_1 = 101;
        if (qp3[102]) n3_1 = 102;
        if (qp2[102]) n2_1 = 102;
        if (qp1[102]) n1_1 = 102;
        if (qp0[102]) n0_1 = 102;
        if (qp3[103]) n3_1 = 103;
        if (qp2[103]) n2_1 = 103;
        if (qp1[103]) n1_1 = 103;
        if (qp0[103]) n0_1 = 103;
        if (qp3[104]) n3_1 = 104;
        if (qp2[104]) n2_1 = 104;
        if (qp1[104]) n1_1 = 104;
        if (qp0[104]) n0_1 = 104;
        if (qp3[105]) n3_1 = 105;
        if (qp2[105]) n2_1 = 105;
        if (qp1[105]) n1_1 = 105;
        if (qp0[105]) n0_1 = 105;
        if (qp3[106]) n3_1 = 106;
        if (qp2[106]) n2_1 = 106;
        if (qp1[106]) n1_1 = 106;
        if (qp0[106]) n0_1 = 106;
        if (qp3[107]) n3_1 = 107;
        if (qp2[107]) n2_1 = 107;
        if (qp1[107]) n1_1 = 107;
        if (qp0[107]) n0_1 = 107;
        if (qp3[108]) n3_1 = 108;
        if (qp2[108]) n2_1 = 108;
        if (qp1[108]) n1_1 = 108;
        if (qp0[108]) n0_1 = 108;
        if (qp3[109]) n3_1 = 109;
        if (qp2[109]) n2_1 = 109;
        if (qp1[109]) n1_1 = 109;
        if (qp0[109]) n0_1 = 109;
        if (qp3[110]) n3_1 = 110;
        if (qp2[110]) n2_1 = 110;
        if (qp1[110]) n1_1 = 110;
        if (qp0[110]) n0_1 = 110;
        if (qp3[111]) n3_1 = 111;
        if (qp2[111]) n2_1 = 111;
        if (qp1[111]) n1_1 = 111;
        if (qp0[111]) n0_1 = 111;
        n3_2 = 7'h7f;
        n2_2 = 7'h7f;
        n1_2 = 7'h7f;
        n0_2 = 7'h7f;
        if (qp3[111]) n3_2 = 111;
        if (qp2[111]) n2_2 = 111;
        if (qp1[111]) n1_2 = 111;
        if (qp0[111]) n0_2 = 111;
        if (qp3[110]) n3_2 = 110;
        if (qp2[110]) n2_2 = 110;
        if (qp1[110]) n1_2 = 110;
        if (qp0[110]) n0_2 = 110;
        if (qp3[109]) n3_2 = 109;
        if (qp2[109]) n2_2 = 109;
        if (qp1[109]) n1_2 = 109;
        if (qp0[109]) n0_2 = 109;
        if (qp3[108]) n3_2 = 108;
        if (qp2[108]) n2_2 = 108;
        if (qp1[108]) n1_2 = 108;
        if (qp0[108]) n0_2 = 108;
        if (qp3[107]) n3_2 = 107;
        if (qp2[107]) n2_2 = 107;
        if (qp1[107]) n1_2 = 107;
        if (qp0[107]) n0_2 = 107;
        if (qp3[106]) n3_2 = 106;
        if (qp2[106]) n2_2 = 106;
        if (qp1[106]) n1_2 = 106;
        if (qp0[106]) n0_2 = 106;
        if (qp3[105]) n3_2 = 105;
        if (qp2[105]) n2_2 = 105;
        if (qp1[105]) n1_2 = 105;
        if (qp0[105]) n0_2 = 105;
        if (qp3[104]) n3_2 = 104;
        if (qp2[104]) n2_2 = 104;
        if (qp1[104]) n1_2 = 104;
        if (qp0[104]) n0_2 = 104;
        if (qp3[103]) n3_2 = 103;
        if (qp2[103]) n2_2 = 103;
        if (qp1[103]) n1_2 = 103;
        if (qp0[103]) n0_2 = 103;
        if (qp3[102]) n3_2 = 102;
        if (qp2[102]) n2_2 = 102;
        if (qp1[102]) n1_2 = 102;
        if (qp0[102]) n0_2 = 102;
        if (qp3[101]) n3_2 = 101;
        if (qp2[101]) n2_2 = 101;
        if (qp1[101]) n1_2 = 101;
        if (qp0[101]) n0_2 = 101;
        if (qp3[100]) n3_2 = 100;
        if (qp2[100]) n2_2 = 100;
        if (qp1[100]) n1_2 = 100;
        if (qp0[100]) n0_2 = 100;
        if (qp3[99]) n3_2 = 99;
        if (qp2[99]) n2_2 = 99;
        if (qp1[99]) n1_2 = 99;
        if (qp0[99]) n0_2 = 99;
        if (qp3[98]) n3_2 = 98;
        if (qp2[98]) n2_2 = 98;
        if (qp1[98]) n1_2 = 98;
        if (qp0[98]) n0_2 = 98;
        if (qp3[97]) n3_2 = 97;
        if (qp2[97]) n2_2 = 97;
        if (qp1[97]) n1_2 = 97;
        if (qp0[97]) n0_2 = 97;
        if (qp3[96]) n3_2 = 96;
        if (qp2[96]) n2_2 = 96;
        if (qp1[96]) n1_2 = 96;
        if (qp0[96]) n0_2 = 96;
        if (qp3[95]) n3_2 = 95;
        if (qp2[95]) n2_2 = 95;
        if (qp1[95]) n1_2 = 95;
        if (qp0[95]) n0_2 = 95;
        if (qp3[94]) n3_2 = 94;
        if (qp2[94]) n2_2 = 94;
        if (qp1[94]) n1_2 = 94;
        if (qp0[94]) n0_2 = 94;
        if (qp3[93]) n3_2 = 93;
        if (qp2[93]) n2_2 = 93;
        if (qp1[93]) n1_2 = 93;
        if (qp0[93]) n0_2 = 93;
        if (qp3[92]) n3_2 = 92;
        if (qp2[92]) n2_2 = 92;
        if (qp1[92]) n1_2 = 92;
        if (qp0[92]) n0_2 = 92;
        if (qp3[91]) n3_2 = 91;
        if (qp2[91]) n2_2 = 91;
        if (qp1[91]) n1_2 = 91;
        if (qp0[91]) n0_2 = 91;
        if (qp3[90]) n3_2 = 90;
        if (qp2[90]) n2_2 = 90;
        if (qp1[90]) n1_2 = 90;
        if (qp0[90]) n0_2 = 90;
        if (qp3[89]) n3_2 = 89;
        if (qp2[89]) n2_2 = 89;
        if (qp1[89]) n1_2 = 89;
        if (qp0[89]) n0_2 = 89;
        if (qp3[88]) n3_2 = 88;
        if (qp2[88]) n2_2 = 88;
        if (qp1[88]) n1_2 = 88;
        if (qp0[88]) n0_2 = 88;
        if (qp3[87]) n3_2 = 87;
        if (qp2[87]) n2_2 = 87;
        if (qp1[87]) n1_2 = 87;
        if (qp0[87]) n0_2 = 87;
        if (qp3[86]) n3_2 = 86;
        if (qp2[86]) n2_2 = 86;
        if (qp1[86]) n1_2 = 86;
        if (qp0[86]) n0_2 = 86;
        if (qp3[85]) n3_2 = 85;
        if (qp2[85]) n2_2 = 85;
        if (qp1[85]) n1_2 = 85;
        if (qp0[85]) n0_2 = 85;
        if (qp3[84]) n3_2 = 84;
        if (qp2[84]) n2_2 = 84;
        if (qp1[84]) n1_2 = 84;
        if (qp0[84]) n0_2 = 84;
        if (qp3[83]) n3_2 = 83;
        if (qp2[83]) n2_2 = 83;
        if (qp1[83]) n1_2 = 83;
        if (qp0[83]) n0_2 = 83;
        if (qp3[82]) n3_2 = 82;
        if (qp2[82]) n2_2 = 82;
        if (qp1[82]) n1_2 = 82;
        if (qp0[82]) n0_2 = 82;
        if (qp3[81]) n3_2 = 81;
        if (qp2[81]) n2_2 = 81;
        if (qp1[81]) n1_2 = 81;
        if (qp0[81]) n0_2 = 81;
        if (qp3[80]) n3_2 = 80;
        if (qp2[80]) n2_2 = 80;
        if (qp1[80]) n1_2 = 80;
        if (qp0[80]) n0_2 = 80;
        if (qp3[79]) n3_2 = 79;
        if (qp2[79]) n2_2 = 79;
        if (qp1[79]) n1_2 = 79;
        if (qp0[79]) n0_2 = 79;
        if (qp3[78]) n3_2 = 78;
        if (qp2[78]) n2_2 = 78;
        if (qp1[78]) n1_2 = 78;
        if (qp0[78]) n0_2 = 78;
        if (qp3[77]) n3_2 = 77;
        if (qp2[77]) n2_2 = 77;
        if (qp1[77]) n1_2 = 77;
        if (qp0[77]) n0_2 = 77;
        if (qp3[76]) n3_2 = 76;
        if (qp2[76]) n2_2 = 76;
        if (qp1[76]) n1_2 = 76;
        if (qp0[76]) n0_2 = 76;
        if (qp3[75]) n3_2 = 75;
        if (qp2[75]) n2_2 = 75;
        if (qp1[75]) n1_2 = 75;
        if (qp0[75]) n0_2 = 75;
        if (qp3[74]) n3_2 = 74;
        if (qp2[74]) n2_2 = 74;
        if (qp1[74]) n1_2 = 74;
        if (qp0[74]) n0_2 = 74;
        if (qp3[73]) n3_2 = 73;
        if (qp2[73]) n2_2 = 73;
        if (qp1[73]) n1_2 = 73;
        if (qp0[73]) n0_2 = 73;
        if (qp3[72]) n3_2 = 72;
        if (qp2[72]) n2_2 = 72;
        if (qp1[72]) n1_2 = 72;
        if (qp0[72]) n0_2 = 72;
        if (qp3[71]) n3_2 = 71;
        if (qp2[71]) n2_2 = 71;
        if (qp1[71]) n1_2 = 71;
        if (qp0[71]) n0_2 = 71;
        if (qp3[70]) n3_2 = 70;
        if (qp2[70]) n2_2 = 70;
        if (qp1[70]) n1_2 = 70;
        if (qp0[70]) n0_2 = 70;
        if (qp3[69]) n3_2 = 69;
        if (qp2[69]) n2_2 = 69;
        if (qp1[69]) n1_2 = 69;
        if (qp0[69]) n0_2 = 69;
        if (qp3[68]) n3_2 = 68;
        if (qp2[68]) n2_2 = 68;
        if (qp1[68]) n1_2 = 68;
        if (qp0[68]) n0_2 = 68;
        if (qp3[67]) n3_2 = 67;
        if (qp2[67]) n2_2 = 67;
        if (qp1[67]) n1_2 = 67;
        if (qp0[67]) n0_2 = 67;
        if (qp3[66]) n3_2 = 66;
        if (qp2[66]) n2_2 = 66;
        if (qp1[66]) n1_2 = 66;
        if (qp0[66]) n0_2 = 66;
        if (qp3[65]) n3_2 = 65;
        if (qp2[65]) n2_2 = 65;
        if (qp1[65]) n1_2 = 65;
        if (qp0[65]) n0_2 = 65;
        if (qp3[64]) n3_2 = 64;
        if (qp2[64]) n2_2 = 64;
        if (qp1[64]) n1_2 = 64;
        if (qp0[64]) n0_2 = 64;
        if (qp3[63]) n3_2 = 63;
        if (qp2[63]) n2_2 = 63;
        if (qp1[63]) n1_2 = 63;
        if (qp0[63]) n0_2 = 63;
        if (qp3[62]) n3_2 = 62;
        if (qp2[62]) n2_2 = 62;
        if (qp1[62]) n1_2 = 62;
        if (qp0[62]) n0_2 = 62;
        if (qp3[61]) n3_2 = 61;
        if (qp2[61]) n2_2 = 61;
        if (qp1[61]) n1_2 = 61;
        if (qp0[61]) n0_2 = 61;
        if (qp3[60]) n3_2 = 60;
        if (qp2[60]) n2_2 = 60;
        if (qp1[60]) n1_2 = 60;
        if (qp0[60]) n0_2 = 60;
        if (qp3[59]) n3_2 = 59;
        if (qp2[59]) n2_2 = 59;
        if (qp1[59]) n1_2 = 59;
        if (qp0[59]) n0_2 = 59;
        if (qp3[58]) n3_2 = 58;
        if (qp2[58]) n2_2 = 58;
        if (qp1[58]) n1_2 = 58;
        if (qp0[58]) n0_2 = 58;
        if (qp3[57]) n3_2 = 57;
        if (qp2[57]) n2_2 = 57;
        if (qp1[57]) n1_2 = 57;
        if (qp0[57]) n0_2 = 57;
        if (qp3[56]) n3_2 = 56;
        if (qp2[56]) n2_2 = 56;
        if (qp1[56]) n1_2 = 56;
        if (qp0[56]) n0_2 = 56;
        if (qp3[55]) n3_2 = 55;
        if (qp2[55]) n2_2 = 55;
        if (qp1[55]) n1_2 = 55;
        if (qp0[55]) n0_2 = 55;
        if (qp3[54]) n3_2 = 54;
        if (qp2[54]) n2_2 = 54;
        if (qp1[54]) n1_2 = 54;
        if (qp0[54]) n0_2 = 54;
        if (qp3[53]) n3_2 = 53;
        if (qp2[53]) n2_2 = 53;
        if (qp1[53]) n1_2 = 53;
        if (qp0[53]) n0_2 = 53;
        if (qp3[52]) n3_2 = 52;
        if (qp2[52]) n2_2 = 52;
        if (qp1[52]) n1_2 = 52;
        if (qp0[52]) n0_2 = 52;
        if (qp3[51]) n3_2 = 51;
        if (qp2[51]) n2_2 = 51;
        if (qp1[51]) n1_2 = 51;
        if (qp0[51]) n0_2 = 51;
        if (qp3[50]) n3_2 = 50;
        if (qp2[50]) n2_2 = 50;
        if (qp1[50]) n1_2 = 50;
        if (qp0[50]) n0_2 = 50;
        if (qp3[49]) n3_2 = 49;
        if (qp2[49]) n2_2 = 49;
        if (qp1[49]) n1_2 = 49;
        if (qp0[49]) n0_2 = 49;
        if (qp3[48]) n3_2 = 48;
        if (qp2[48]) n2_2 = 48;
        if (qp1[48]) n1_2 = 48;
        if (qp0[48]) n0_2 = 48;
        if (qp3[47]) n3_2 = 47;
        if (qp2[47]) n2_2 = 47;
        if (qp1[47]) n1_2 = 47;
        if (qp0[47]) n0_2 = 47;
        if (qp3[46]) n3_2 = 46;
        if (qp2[46]) n2_2 = 46;
        if (qp1[46]) n1_2 = 46;
        if (qp0[46]) n0_2 = 46;
        if (qp3[45]) n3_2 = 45;
        if (qp2[45]) n2_2 = 45;
        if (qp1[45]) n1_2 = 45;
        if (qp0[45]) n0_2 = 45;
        if (qp3[44]) n3_2 = 44;
        if (qp2[44]) n2_2 = 44;
        if (qp1[44]) n1_2 = 44;
        if (qp0[44]) n0_2 = 44;
        if (qp3[43]) n3_2 = 43;
        if (qp2[43]) n2_2 = 43;
        if (qp1[43]) n1_2 = 43;
        if (qp0[43]) n0_2 = 43;
        if (qp3[42]) n3_2 = 42;
        if (qp2[42]) n2_2 = 42;
        if (qp1[42]) n1_2 = 42;
        if (qp0[42]) n0_2 = 42;
        if (qp3[41]) n3_2 = 41;
        if (qp2[41]) n2_2 = 41;
        if (qp1[41]) n1_2 = 41;
        if (qp0[41]) n0_2 = 41;
        if (qp3[40]) n3_2 = 40;
        if (qp2[40]) n2_2 = 40;
        if (qp1[40]) n1_2 = 40;
        if (qp0[40]) n0_2 = 40;
        if (qp3[39]) n3_2 = 39;
        if (qp2[39]) n2_2 = 39;
        if (qp1[39]) n1_2 = 39;
        if (qp0[39]) n0_2 = 39;
        if (qp3[38]) n3_2 = 38;
        if (qp2[38]) n2_2 = 38;
        if (qp1[38]) n1_2 = 38;
        if (qp0[38]) n0_2 = 38;
        if (qp3[37]) n3_2 = 37;
        if (qp2[37]) n2_2 = 37;
        if (qp1[37]) n1_2 = 37;
        if (qp0[37]) n0_2 = 37;
        if (qp3[36]) n3_2 = 36;
        if (qp2[36]) n2_2 = 36;
        if (qp1[36]) n1_2 = 36;
        if (qp0[36]) n0_2 = 36;
        if (qp3[35]) n3_2 = 35;
        if (qp2[35]) n2_2 = 35;
        if (qp1[35]) n1_2 = 35;
        if (qp0[35]) n0_2 = 35;
        if (qp3[34]) n3_2 = 34;
        if (qp2[34]) n2_2 = 34;
        if (qp1[34]) n1_2 = 34;
        if (qp0[34]) n0_2 = 34;
        if (qp3[33]) n3_2 = 33;
        if (qp2[33]) n2_2 = 33;
        if (qp1[33]) n1_2 = 33;
        if (qp0[33]) n0_2 = 33;
        if (qp3[32]) n3_2 = 32;
        if (qp2[32]) n2_2 = 32;
        if (qp1[32]) n1_2 = 32;
        if (qp0[32]) n0_2 = 32;
        if (qp3[31]) n3_2 = 31;
        if (qp2[31]) n2_2 = 31;
        if (qp1[31]) n1_2 = 31;
        if (qp0[31]) n0_2 = 31;
        if (qp3[30]) n3_2 = 30;
        if (qp2[30]) n2_2 = 30;
        if (qp1[30]) n1_2 = 30;
        if (qp0[30]) n0_2 = 30;
        if (qp3[29]) n3_2 = 29;
        if (qp2[29]) n2_2 = 29;
        if (qp1[29]) n1_2 = 29;
        if (qp0[29]) n0_2 = 29;
        if (qp3[28]) n3_2 = 28;
        if (qp2[28]) n2_2 = 28;
        if (qp1[28]) n1_2 = 28;
        if (qp0[28]) n0_2 = 28;
        if (qp3[27]) n3_2 = 27;
        if (qp2[27]) n2_2 = 27;
        if (qp1[27]) n1_2 = 27;
        if (qp0[27]) n0_2 = 27;
        if (qp3[26]) n3_2 = 26;
        if (qp2[26]) n2_2 = 26;
        if (qp1[26]) n1_2 = 26;
        if (qp0[26]) n0_2 = 26;
        if (qp3[25]) n3_2 = 25;
        if (qp2[25]) n2_2 = 25;
        if (qp1[25]) n1_2 = 25;
        if (qp0[25]) n0_2 = 25;
        if (qp3[24]) n3_2 = 24;
        if (qp2[24]) n2_2 = 24;
        if (qp1[24]) n1_2 = 24;
        if (qp0[24]) n0_2 = 24;
        if (qp3[23]) n3_2 = 23;
        if (qp2[23]) n2_2 = 23;
        if (qp1[23]) n1_2 = 23;
        if (qp0[23]) n0_2 = 23;
        if (qp3[22]) n3_2 = 22;
        if (qp2[22]) n2_2 = 22;
        if (qp1[22]) n1_2 = 22;
        if (qp0[22]) n0_2 = 22;
        if (qp3[21]) n3_2 = 21;
        if (qp2[21]) n2_2 = 21;
        if (qp1[21]) n1_2 = 21;
        if (qp0[21]) n0_2 = 21;
        if (qp3[20]) n3_2 = 20;
        if (qp2[20]) n2_2 = 20;
        if (qp1[20]) n1_2 = 20;
        if (qp0[20]) n0_2 = 20;
        if (qp3[19]) n3_2 = 19;
        if (qp2[19]) n2_2 = 19;
        if (qp1[19]) n1_2 = 19;
        if (qp0[19]) n0_2 = 19;
        if (qp3[18]) n3_2 = 18;
        if (qp2[18]) n2_2 = 18;
        if (qp1[18]) n1_2 = 18;
        if (qp0[18]) n0_2 = 18;
        if (qp3[17]) n3_2 = 17;
        if (qp2[17]) n2_2 = 17;
        if (qp1[17]) n1_2 = 17;
        if (qp0[17]) n0_2 = 17;
        if (qp3[16]) n3_2 = 16;
        if (qp2[16]) n2_2 = 16;
        if (qp1[16]) n1_2 = 16;
        if (qp0[16]) n0_2 = 16;
        if (qp3[15]) n3_2 = 15;
        if (qp2[15]) n2_2 = 15;
        if (qp1[15]) n1_2 = 15;
        if (qp0[15]) n0_2 = 15;
        if (qp3[14]) n3_2 = 14;
        if (qp2[14]) n2_2 = 14;
        if (qp1[14]) n1_2 = 14;
        if (qp0[14]) n0_2 = 14;
        if (qp3[13]) n3_2 = 13;
        if (qp2[13]) n2_2 = 13;
        if (qp1[13]) n1_2 = 13;
        if (qp0[13]) n0_2 = 13;
        if (qp3[12]) n3_2 = 12;
        if (qp2[12]) n2_2 = 12;
        if (qp1[12]) n1_2 = 12;
        if (qp0[12]) n0_2 = 12;
        if (qp3[11]) n3_2 = 11;
        if (qp2[11]) n2_2 = 11;
        if (qp1[11]) n1_2 = 11;
        if (qp0[11]) n0_2 = 11;
        if (qp3[10]) n3_2 = 10;
        if (qp2[10]) n2_2 = 10;
        if (qp1[10]) n1_2 = 10;
        if (qp0[10]) n0_2 = 10;
        if (qp3[9]) n3_2 = 9;
        if (qp2[9]) n2_2 = 9;
        if (qp1[9]) n1_2 = 9;
        if (qp0[9]) n0_2 = 9;
        if (qp3[8]) n3_2 = 8;
        if (qp2[8]) n2_2 = 8;
        if (qp1[8]) n1_2 = 8;
        if (qp0[8]) n0_2 = 8;
        if (qp3[7]) n3_2 = 7;
        if (qp2[7]) n2_2 = 7;
        if (qp1[7]) n1_2 = 7;
        if (qp0[7]) n0_2 = 7;
        if (qp3[6]) n3_2 = 6;
        if (qp2[6]) n2_2 = 6;
        if (qp1[6]) n1_2 = 6;
        if (qp0[6]) n0_2 = 6;
        if (qp3[5]) n3_2 = 5;
        if (qp2[5]) n2_2 = 5;
        if (qp1[5]) n1_2 = 5;
        if (qp0[5]) n0_2 = 5;
        if (qp3[4]) n3_2 = 4;
        if (qp2[4]) n2_2 = 4;
        if (qp1[4]) n1_2 = 4;
        if (qp0[4]) n0_2 = 4;
        if (qp3[3]) n3_2 = 3;
        if (qp2[3]) n2_2 = 3;
        if (qp1[3]) n1_2 = 3;
        if (qp0[3]) n0_2 = 3;
        if (qp3[2]) n3_2 = 2;
        if (qp2[2]) n2_2 = 2;
        if (qp1[2]) n1_2 = 2;
        if (qp0[2]) n0_2 = 2;
        if (qp3[1]) n3_2 = 1;
        if (qp2[1]) n2_2 = 1;
        if (qp1[1]) n1_2 = 1;
        if (qp0[1]) n0_2 = 1;
        if (qp3[0]) n3_2 = 0;
        if (qp2[0]) n2_2 = 0;
        if (qp1[0]) n1_2 = 0;
        if (qp0[0]) n0_2 = 0;
        q1 = 0;
        q2 = 0;
        w1 = 0;
        w2 = 0;
        v1 = 0;
        v2 = 0;
        if (n3_1 != 7'h7f) 
        begin
            w1 = n3_1;
            q1 = 3;
            v1 = 1;
            if (n3_1 != n3_2) 
            begin
                w2 = n3_2;
                q2 = 3;
                v2 = 1;
            end
            else if (n2_1 != 7'h7f) 
            begin
                w2 = n2_1;
                q2 = 2;
                v2 = 1;
            end
            else if (n1_1 != 7'h7f) 
            begin
                w2 = n1_1;
                q2 = 1;
                v2 = 1;
            end
            else if (n0_1 != 7'h7f) 
            begin
                w2 = n0_1;
                q2 = 0;
                v2 = 1;
            end
        end
        else 
        begin
            if (n2_1 != 7'h7f) 
            begin
                w1 = n2_1;
                q1 = 2;
                v1 = 1;
                if (n2_1 != n2_2) 
                begin
                    w2 = n2_2;
                    q2 = 2;
                    v2 = 1;
                end
                else if (n1_1 != 7'h7f) 
                begin
                    w2 = n1_1;
                    q2 = 1;
                    v2 = 1;
                end
                else if (n0_1 != 7'h7f) 
                begin
                    w2 = n0_1;
                    q2 = 0;
                    v2 = 1;
                end
            end
            else 
            begin
                if (n1_1 != 7'h7f) 
                begin
                    w1 = n1_1;
                    q1 = 1;
                    v1 = 1;
                    if (n1_1 != n1_2) 
                    begin
                        w2 = n1_2;
                        q2 = 1;
                        v2 = 1;
                    end
                    else if (n0_1 != 7'h7f) 
                    begin
                        w2 = n0_1;
                        q2 = 0;
                        v2 = 1;
                    end
                end
                else 
                begin
                    if (n0_1 != 7'h7f) 
                    begin
                        w1 = n0_1;
                        q1 = 0;
                        v1 = 1;
                        if (n0_1 != n0_2) 
                        begin
                            w2 = n0_2;
                            q2 = 0;
                            v2 = 1;
                        end
                    end
                end
            end
        end
    end
endmodule
